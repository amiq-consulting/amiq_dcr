/******************************************************************************
 * (C) Copyright 2015 AMIQ Consulting
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * NAME:        amiq_dcr_ex_ms_defines.sv
 * PROJECT:     amiq_dcr
 * Description: This file contains the declaration of all the used defines
 *******************************************************************************/

`ifndef AMIQ_DCR_EX_MS_DEFINES_SV
	//protection against multiple includes
	`define AMIQ_DCR_EX_MS_DEFINES_SV

	//number of registers
	`define AMIQ_DCR_EX_MS_NUMBER_OF_REGS 32

`endif

